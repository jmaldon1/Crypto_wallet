// crypto_wallet2_nios_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module crypto_wallet2_nios_tb (
	);

	wire         crypto_wallet2_nios_inst_clk_bfm_clk_clk;                                  // crypto_wallet2_nios_inst_clk_bfm:clk -> [crypto_wallet2_nios_inst:clk_clk, crypto_wallet2_nios_inst_reset_bfm:clk]
	wire         crypto_wallet2_nios_inst_epcs_flash_controller_external_dclk;              // crypto_wallet2_nios_inst:epcs_flash_controller_external_dclk -> crypto_wallet2_nios_inst_epcs_flash_controller_external_bfm:sig_dclk
	wire         crypto_wallet2_nios_inst_epcs_flash_controller_external_sce;               // crypto_wallet2_nios_inst:epcs_flash_controller_external_sce -> crypto_wallet2_nios_inst_epcs_flash_controller_external_bfm:sig_sce
	wire   [0:0] crypto_wallet2_nios_inst_epcs_flash_controller_external_bfm_conduit_data0; // crypto_wallet2_nios_inst_epcs_flash_controller_external_bfm:sig_data0 -> crypto_wallet2_nios_inst:epcs_flash_controller_external_data0
	wire         crypto_wallet2_nios_inst_epcs_flash_controller_external_sdo;               // crypto_wallet2_nios_inst:epcs_flash_controller_external_sdo -> crypto_wallet2_nios_inst_epcs_flash_controller_external_bfm:sig_sdo
	wire   [7:0] crypto_wallet2_nios_inst_po_led_external_connection_export;                // crypto_wallet2_nios_inst:po_led_external_connection_export -> crypto_wallet2_nios_inst_po_led_external_connection_bfm:sig_export
	wire         crypto_wallet2_nios_inst_sdram_wire_cs_n;                                  // crypto_wallet2_nios_inst:sdram_wire_cs_n -> crypto_wallet2_nios_inst_sdram_wire_bfm:sig_cs_n
	wire   [1:0] crypto_wallet2_nios_inst_sdram_wire_dqm;                                   // crypto_wallet2_nios_inst:sdram_wire_dqm -> crypto_wallet2_nios_inst_sdram_wire_bfm:sig_dqm
	wire         crypto_wallet2_nios_inst_sdram_wire_cas_n;                                 // crypto_wallet2_nios_inst:sdram_wire_cas_n -> crypto_wallet2_nios_inst_sdram_wire_bfm:sig_cas_n
	wire         crypto_wallet2_nios_inst_sdram_wire_ras_n;                                 // crypto_wallet2_nios_inst:sdram_wire_ras_n -> crypto_wallet2_nios_inst_sdram_wire_bfm:sig_ras_n
	wire         crypto_wallet2_nios_inst_sdram_wire_we_n;                                  // crypto_wallet2_nios_inst:sdram_wire_we_n -> crypto_wallet2_nios_inst_sdram_wire_bfm:sig_we_n
	wire  [12:0] crypto_wallet2_nios_inst_sdram_wire_addr;                                  // crypto_wallet2_nios_inst:sdram_wire_addr -> crypto_wallet2_nios_inst_sdram_wire_bfm:sig_addr
	wire         crypto_wallet2_nios_inst_sdram_wire_cke;                                   // crypto_wallet2_nios_inst:sdram_wire_cke -> crypto_wallet2_nios_inst_sdram_wire_bfm:sig_cke
	wire  [15:0] crypto_wallet2_nios_inst_sdram_wire_dq;                                    // [] -> [crypto_wallet2_nios_inst:sdram_wire_dq, crypto_wallet2_nios_inst_sdram_wire_bfm:sig_dq]
	wire   [1:0] crypto_wallet2_nios_inst_sdram_wire_ba;                                    // crypto_wallet2_nios_inst:sdram_wire_ba -> crypto_wallet2_nios_inst_sdram_wire_bfm:sig_ba
	wire         crypto_wallet2_nios_inst_uart_external_connection_txd;                     // crypto_wallet2_nios_inst:uart_external_connection_txd -> crypto_wallet2_nios_inst_uart_external_connection_bfm:sig_txd
	wire   [0:0] crypto_wallet2_nios_inst_uart_external_connection_bfm_conduit_rxd;         // crypto_wallet2_nios_inst_uart_external_connection_bfm:sig_rxd -> crypto_wallet2_nios_inst:uart_external_connection_rxd
	wire         crypto_wallet2_nios_inst_reset_bfm_reset_reset;                            // crypto_wallet2_nios_inst_reset_bfm:reset -> crypto_wallet2_nios_inst:reset_reset_n

	crypto_wallet2_nios crypto_wallet2_nios_inst (
		.clk_clk                              (crypto_wallet2_nios_inst_clk_bfm_clk_clk),                                  //                            clk.clk
		.epcs_flash_controller_external_dclk  (crypto_wallet2_nios_inst_epcs_flash_controller_external_dclk),              // epcs_flash_controller_external.dclk
		.epcs_flash_controller_external_sce   (crypto_wallet2_nios_inst_epcs_flash_controller_external_sce),               //                               .sce
		.epcs_flash_controller_external_sdo   (crypto_wallet2_nios_inst_epcs_flash_controller_external_sdo),               //                               .sdo
		.epcs_flash_controller_external_data0 (crypto_wallet2_nios_inst_epcs_flash_controller_external_bfm_conduit_data0), //                               .data0
		.po_led_external_connection_export    (crypto_wallet2_nios_inst_po_led_external_connection_export),                //     po_led_external_connection.export
		.reset_reset_n                        (crypto_wallet2_nios_inst_reset_bfm_reset_reset),                            //                          reset.reset_n
		.sdram_wire_addr                      (crypto_wallet2_nios_inst_sdram_wire_addr),                                  //                     sdram_wire.addr
		.sdram_wire_ba                        (crypto_wallet2_nios_inst_sdram_wire_ba),                                    //                               .ba
		.sdram_wire_cas_n                     (crypto_wallet2_nios_inst_sdram_wire_cas_n),                                 //                               .cas_n
		.sdram_wire_cke                       (crypto_wallet2_nios_inst_sdram_wire_cke),                                   //                               .cke
		.sdram_wire_cs_n                      (crypto_wallet2_nios_inst_sdram_wire_cs_n),                                  //                               .cs_n
		.sdram_wire_dq                        (crypto_wallet2_nios_inst_sdram_wire_dq),                                    //                               .dq
		.sdram_wire_dqm                       (crypto_wallet2_nios_inst_sdram_wire_dqm),                                   //                               .dqm
		.sdram_wire_ras_n                     (crypto_wallet2_nios_inst_sdram_wire_ras_n),                                 //                               .ras_n
		.sdram_wire_we_n                      (crypto_wallet2_nios_inst_sdram_wire_we_n),                                  //                               .we_n
		.uart_external_connection_rxd         (crypto_wallet2_nios_inst_uart_external_connection_bfm_conduit_rxd),         //       uart_external_connection.rxd
		.uart_external_connection_txd         (crypto_wallet2_nios_inst_uart_external_connection_txd)                      //                               .txd
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) crypto_wallet2_nios_inst_clk_bfm (
		.clk (crypto_wallet2_nios_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm crypto_wallet2_nios_inst_epcs_flash_controller_external_bfm (
		.sig_data0 (crypto_wallet2_nios_inst_epcs_flash_controller_external_bfm_conduit_data0), // conduit.data0
		.sig_dclk  (crypto_wallet2_nios_inst_epcs_flash_controller_external_dclk),              //        .dclk
		.sig_sce   (crypto_wallet2_nios_inst_epcs_flash_controller_external_sce),               //        .sce
		.sig_sdo   (crypto_wallet2_nios_inst_epcs_flash_controller_external_sdo)                //        .sdo
	);

	altera_conduit_bfm_0002 crypto_wallet2_nios_inst_po_led_external_connection_bfm (
		.sig_export (crypto_wallet2_nios_inst_po_led_external_connection_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) crypto_wallet2_nios_inst_reset_bfm (
		.reset (crypto_wallet2_nios_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (crypto_wallet2_nios_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0003 crypto_wallet2_nios_inst_sdram_wire_bfm (
		.sig_addr  (crypto_wallet2_nios_inst_sdram_wire_addr),  // conduit.addr
		.sig_ba    (crypto_wallet2_nios_inst_sdram_wire_ba),    //        .ba
		.sig_cas_n (crypto_wallet2_nios_inst_sdram_wire_cas_n), //        .cas_n
		.sig_cke   (crypto_wallet2_nios_inst_sdram_wire_cke),   //        .cke
		.sig_cs_n  (crypto_wallet2_nios_inst_sdram_wire_cs_n),  //        .cs_n
		.sig_dq    (crypto_wallet2_nios_inst_sdram_wire_dq),    //        .dq
		.sig_dqm   (crypto_wallet2_nios_inst_sdram_wire_dqm),   //        .dqm
		.sig_ras_n (crypto_wallet2_nios_inst_sdram_wire_ras_n), //        .ras_n
		.sig_we_n  (crypto_wallet2_nios_inst_sdram_wire_we_n)   //        .we_n
	);

	altera_conduit_bfm_0004 crypto_wallet2_nios_inst_uart_external_connection_bfm (
		.sig_rxd (crypto_wallet2_nios_inst_uart_external_connection_bfm_conduit_rxd), // conduit.rxd
		.sig_txd (crypto_wallet2_nios_inst_uart_external_connection_txd)              //        .txd
	);

endmodule
