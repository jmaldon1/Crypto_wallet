-- crypto_wallet.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity crypto_wallet is
	port (
		clk_clk                                     : in    std_logic                     := '0';             --                                  clk.clk
		epcs_flash_controller_dclk                  : out   std_logic;                                        --                epcs_flash_controller.dclk
		epcs_flash_controller_sce                   : out   std_logic;                                        --                                     .sce
		epcs_flash_controller_sdo                   : out   std_logic;                                        --                                     .sdo
		epcs_flash_controller_data0                 : in    std_logic                     := '0';             --                                     .data0
		pi_gpio0_external_connection_export         : in    std_logic_vector(1 downto 0)  := (others => '0'); --         pi_gpio0_external_connection.export
		pi_gpio1_external_connection_export         : in    std_logic_vector(1 downto 0)  := (others => '0'); --         pi_gpio1_external_connection.export
		pi_gpio2_external_connection_export         : in    std_logic_vector(2 downto 0)  := (others => '0'); --         pi_gpio2_external_connection.export
		pi_key_external_connection_export           : in    std_logic_vector(1 downto 0)  := (others => '0'); --           pi_key_external_connection.export
		pi_sw_external_connection_export            : in    std_logic_vector(3 downto 0)  := (others => '0'); --            pi_sw_external_connection.export
		pio_gpio0_33to32_external_connection_export : inout std_logic_vector(1 downto 0)  := (others => '0'); -- pio_gpio0_33to32_external_connection.export
		pio_gpio0_external_connection_export        : inout std_logic_vector(31 downto 0) := (others => '0'); --        pio_gpio0_external_connection.export
		pio_gpio1_33to32_external_connection_export : inout std_logic_vector(1 downto 0)  := (others => '0'); -- pio_gpio1_33to32_external_connection.export
		pio_gpio1_external_connection_export        : inout std_logic_vector(31 downto 0) := (others => '0'); --        pio_gpio1_external_connection.export
		pio_gpio2_external_connection_export        : inout std_logic_vector(12 downto 0) := (others => '0'); --        pio_gpio2_external_connection.export
		po_led_external_connection_export           : out   std_logic_vector(7 downto 0);                     --           po_led_external_connection.export
		reset_n_reset_n                             : in    std_logic                     := '0';             --                              reset_n.reset_n
		sdram_addr                                  : out   std_logic_vector(12 downto 0);                    --                                sdram.addr
		sdram_ba                                    : out   std_logic_vector(1 downto 0);                     --                                     .ba
		sdram_cas_n                                 : out   std_logic;                                        --                                     .cas_n
		sdram_cke                                   : out   std_logic;                                        --                                     .cke
		sdram_cs_n                                  : out   std_logic;                                        --                                     .cs_n
		sdram_dq                                    : inout std_logic_vector(15 downto 0) := (others => '0'); --                                     .dq
		sdram_dqm                                   : out   std_logic_vector(1 downto 0);                     --                                     .dqm
		sdram_ras_n                                 : out   std_logic;                                        --                                     .ras_n
		sdram_we_n                                  : out   std_logic                                         --                                     .we_n
	);
end entity crypto_wallet;

architecture rtl of crypto_wallet is
	component crypto_wallet_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(25 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component crypto_wallet_cpu;

	component crypto_wallet_epcs_flash_controller is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read_n     : in  std_logic                     := 'X';             -- read_n
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq        : out std_logic;                                        -- irq
			dclk       : out std_logic;                                        -- export
			sce        : out std_logic;                                        -- export
			sdo        : out std_logic;                                        -- export
			data0      : in  std_logic                     := 'X'              -- export
		);
	end component crypto_wallet_epcs_flash_controller;

	component crypto_wallet_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component crypto_wallet_jtag_uart;

	component crypto_wallet_onchip_memory2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component crypto_wallet_onchip_memory2;

	component crypto_wallet_pi_gpio0 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component crypto_wallet_pi_gpio0;

	component crypto_wallet_pi_gpio2 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- export
		);
	end component crypto_wallet_pi_gpio2;

	component crypto_wallet_pi_sw is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component crypto_wallet_pi_sw;

	component crypto_wallet_pio_gpio0_31to0 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component crypto_wallet_pio_gpio0_31to0;

	component crypto_wallet_pio_gpio0_33to32 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component crypto_wallet_pio_gpio0_33to32;

	component crypto_wallet_pio_gpio2 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(12 downto 0) := (others => 'X')  -- export
		);
	end component crypto_wallet_pio_gpio2;

	component crypto_wallet_po_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component crypto_wallet_po_led;

	component crypto_wallet_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component crypto_wallet_sdram;

	component crypto_wallet_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component crypto_wallet_sysid;

	component crypto_wallet_mm_interconnect_0 is
		port (
			clk_50_clk_clk                                     : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                            : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                        : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                               : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                              : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                        : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                     : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                 : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                        : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_debug_mem_slave_address                        : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                          : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                           : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                    : out std_logic;                                        -- debugaccess
			epcs_flash_controller_epcs_control_port_address    : out std_logic_vector(8 downto 0);                     -- address
			epcs_flash_controller_epcs_control_port_write      : out std_logic;                                        -- write
			epcs_flash_controller_epcs_control_port_read       : out std_logic;                                        -- read
			epcs_flash_controller_epcs_control_port_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			epcs_flash_controller_epcs_control_port_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			epcs_flash_controller_epcs_control_port_chipselect : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                  : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                   : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect             : out std_logic;                                        -- chipselect
			onchip_memory2_s1_address                          : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_s1_write                            : out std_logic;                                        -- write
			onchip_memory2_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_s1_chipselect                       : out std_logic;                                        -- chipselect
			onchip_memory2_s1_clken                            : out std_logic;                                        -- clken
			pi_gpio0_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			pi_gpio0_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pi_gpio1_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			pi_gpio1_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pi_gpio2_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			pi_gpio2_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pi_key_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			pi_key_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pi_sw_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			pi_sw_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_gpio0_31to0_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			pio_gpio0_31to0_s1_write                           : out std_logic;                                        -- write
			pio_gpio0_31to0_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_gpio0_31to0_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			pio_gpio0_31to0_s1_chipselect                      : out std_logic;                                        -- chipselect
			pio_gpio0_33to32_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			pio_gpio0_33to32_s1_write                          : out std_logic;                                        -- write
			pio_gpio0_33to32_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_gpio0_33to32_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			pio_gpio0_33to32_s1_chipselect                     : out std_logic;                                        -- chipselect
			pio_gpio1_31to0_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			pio_gpio1_31to0_s1_write                           : out std_logic;                                        -- write
			pio_gpio1_31to0_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_gpio1_31to0_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			pio_gpio1_31to0_s1_chipselect                      : out std_logic;                                        -- chipselect
			pio_gpio1_33to32_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			pio_gpio1_33to32_s1_write                          : out std_logic;                                        -- write
			pio_gpio1_33to32_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_gpio1_33to32_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			pio_gpio1_33to32_s1_chipselect                     : out std_logic;                                        -- chipselect
			pio_gpio2_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pio_gpio2_s1_write                                 : out std_logic;                                        -- write
			pio_gpio2_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_gpio2_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pio_gpio2_s1_chipselect                            : out std_logic;                                        -- chipselect
			po_led_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			po_led_s1_write                                    : out std_logic;                                        -- write
			po_led_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			po_led_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			po_led_s1_chipselect                               : out std_logic;                                        -- chipselect
			sdram_s1_address                                   : out std_logic_vector(23 downto 0);                    -- address
			sdram_s1_write                                     : out std_logic;                                        -- write
			sdram_s1_read                                      : out std_logic;                                        -- read
			sdram_s1_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                             : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                : out std_logic;                                        -- chipselect
			sysid_control_slave_address                        : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component crypto_wallet_mm_interconnect_0;

	component crypto_wallet_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component crypto_wallet_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_data_master_readdata                                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                               : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                               : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                   : std_logic_vector(25 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                                : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                      : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                                     : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                                 : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                            : std_logic_vector(25 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                               : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect                  : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                    : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest                 : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                        : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                       : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                            : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                            : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                         : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                         : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                                : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                               : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect      : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_chipselect -> epcs_flash_controller:chipselect
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata        : std_logic_vector(31 downto 0); -- epcs_flash_controller:readdata -> mm_interconnect_0:epcs_flash_controller_epcs_control_port_readdata
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_address -> epcs_flash_controller:address
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_read            : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_read -> mm_interconnect_0_epcs_flash_controller_epcs_control_port_read:in
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_write           : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_write -> mm_interconnect_0_epcs_flash_controller_epcs_control_port_write:in
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_writedata -> epcs_flash_controller:writedata
	signal mm_interconnect_0_po_led_s1_chipselect                                    : std_logic;                     -- mm_interconnect_0:po_led_s1_chipselect -> po_led:chipselect
	signal mm_interconnect_0_po_led_s1_readdata                                      : std_logic_vector(31 downto 0); -- po_led:readdata -> mm_interconnect_0:po_led_s1_readdata
	signal mm_interconnect_0_po_led_s1_address                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:po_led_s1_address -> po_led:address
	signal mm_interconnect_0_po_led_s1_write                                         : std_logic;                     -- mm_interconnect_0:po_led_s1_write -> mm_interconnect_0_po_led_s1_write:in
	signal mm_interconnect_0_po_led_s1_writedata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:po_led_s1_writedata -> po_led:writedata
	signal mm_interconnect_0_onchip_memory2_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	signal mm_interconnect_0_onchip_memory2_s1_readdata                              : std_logic_vector(31 downto 0); -- onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	signal mm_interconnect_0_onchip_memory2_s1_address                               : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	signal mm_interconnect_0_onchip_memory2_s1_byteenable                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	signal mm_interconnect_0_onchip_memory2_s1_write                                 : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	signal mm_interconnect_0_onchip_memory2_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	signal mm_interconnect_0_onchip_memory2_s1_clken                                 : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	signal mm_interconnect_0_pi_key_s1_readdata                                      : std_logic_vector(31 downto 0); -- pi_key:readdata -> mm_interconnect_0:pi_key_s1_readdata
	signal mm_interconnect_0_pi_key_s1_address                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pi_key_s1_address -> pi_key:address
	signal mm_interconnect_0_pi_sw_s1_readdata                                       : std_logic_vector(31 downto 0); -- pi_sw:readdata -> mm_interconnect_0:pi_sw_s1_readdata
	signal mm_interconnect_0_pi_sw_s1_address                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pi_sw_s1_address -> pi_sw:address
	signal mm_interconnect_0_sdram_s1_chipselect                                     : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                       : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                    : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                        : std_logic_vector(23 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                           : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                                  : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                          : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_pi_gpio1_s1_readdata                                    : std_logic_vector(31 downto 0); -- pi_gpio1:readdata -> mm_interconnect_0:pi_gpio1_s1_readdata
	signal mm_interconnect_0_pi_gpio1_s1_address                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pi_gpio1_s1_address -> pi_gpio1:address
	signal mm_interconnect_0_pi_gpio0_s1_readdata                                    : std_logic_vector(31 downto 0); -- pi_gpio0:readdata -> mm_interconnect_0:pi_gpio0_s1_readdata
	signal mm_interconnect_0_pi_gpio0_s1_address                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pi_gpio0_s1_address -> pi_gpio0:address
	signal mm_interconnect_0_pi_gpio2_s1_readdata                                    : std_logic_vector(31 downto 0); -- pi_gpio2:readdata -> mm_interconnect_0:pi_gpio2_s1_readdata
	signal mm_interconnect_0_pi_gpio2_s1_address                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pi_gpio2_s1_address -> pi_gpio2:address
	signal mm_interconnect_0_pio_gpio2_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:pio_gpio2_s1_chipselect -> pio_gpio2:chipselect
	signal mm_interconnect_0_pio_gpio2_s1_readdata                                   : std_logic_vector(31 downto 0); -- pio_gpio2:readdata -> mm_interconnect_0:pio_gpio2_s1_readdata
	signal mm_interconnect_0_pio_gpio2_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_gpio2_s1_address -> pio_gpio2:address
	signal mm_interconnect_0_pio_gpio2_s1_write                                      : std_logic;                     -- mm_interconnect_0:pio_gpio2_s1_write -> mm_interconnect_0_pio_gpio2_s1_write:in
	signal mm_interconnect_0_pio_gpio2_s1_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_gpio2_s1_writedata -> pio_gpio2:writedata
	signal mm_interconnect_0_pio_gpio0_31to0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:pio_gpio0_31to0_s1_chipselect -> pio_gpio0_31to0:chipselect
	signal mm_interconnect_0_pio_gpio0_31to0_s1_readdata                             : std_logic_vector(31 downto 0); -- pio_gpio0_31to0:readdata -> mm_interconnect_0:pio_gpio0_31to0_s1_readdata
	signal mm_interconnect_0_pio_gpio0_31to0_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_gpio0_31to0_s1_address -> pio_gpio0_31to0:address
	signal mm_interconnect_0_pio_gpio0_31to0_s1_write                                : std_logic;                     -- mm_interconnect_0:pio_gpio0_31to0_s1_write -> mm_interconnect_0_pio_gpio0_31to0_s1_write:in
	signal mm_interconnect_0_pio_gpio0_31to0_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_gpio0_31to0_s1_writedata -> pio_gpio0_31to0:writedata
	signal mm_interconnect_0_pio_gpio1_31to0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:pio_gpio1_31to0_s1_chipselect -> pio_gpio1_31to0:chipselect
	signal mm_interconnect_0_pio_gpio1_31to0_s1_readdata                             : std_logic_vector(31 downto 0); -- pio_gpio1_31to0:readdata -> mm_interconnect_0:pio_gpio1_31to0_s1_readdata
	signal mm_interconnect_0_pio_gpio1_31to0_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_gpio1_31to0_s1_address -> pio_gpio1_31to0:address
	signal mm_interconnect_0_pio_gpio1_31to0_s1_write                                : std_logic;                     -- mm_interconnect_0:pio_gpio1_31to0_s1_write -> mm_interconnect_0_pio_gpio1_31to0_s1_write:in
	signal mm_interconnect_0_pio_gpio1_31to0_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_gpio1_31to0_s1_writedata -> pio_gpio1_31to0:writedata
	signal mm_interconnect_0_pio_gpio0_33to32_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:pio_gpio0_33to32_s1_chipselect -> pio_gpio0_33to32:chipselect
	signal mm_interconnect_0_pio_gpio0_33to32_s1_readdata                            : std_logic_vector(31 downto 0); -- pio_gpio0_33to32:readdata -> mm_interconnect_0:pio_gpio0_33to32_s1_readdata
	signal mm_interconnect_0_pio_gpio0_33to32_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_gpio0_33to32_s1_address -> pio_gpio0_33to32:address
	signal mm_interconnect_0_pio_gpio0_33to32_s1_write                               : std_logic;                     -- mm_interconnect_0:pio_gpio0_33to32_s1_write -> mm_interconnect_0_pio_gpio0_33to32_s1_write:in
	signal mm_interconnect_0_pio_gpio0_33to32_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_gpio0_33to32_s1_writedata -> pio_gpio0_33to32:writedata
	signal mm_interconnect_0_pio_gpio1_33to32_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:pio_gpio1_33to32_s1_chipselect -> pio_gpio1_33to32:chipselect
	signal mm_interconnect_0_pio_gpio1_33to32_s1_readdata                            : std_logic_vector(31 downto 0); -- pio_gpio1_33to32:readdata -> mm_interconnect_0:pio_gpio1_33to32_s1_readdata
	signal mm_interconnect_0_pio_gpio1_33to32_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_gpio1_33to32_s1_address -> pio_gpio1_33to32:address
	signal mm_interconnect_0_pio_gpio1_33to32_s1_write                               : std_logic;                     -- mm_interconnect_0:pio_gpio1_33to32_s1_write -> mm_interconnect_0_pio_gpio1_33to32_s1_write:in
	signal mm_interconnect_0_pio_gpio1_33to32_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_gpio1_33to32_s1_writedata -> pio_gpio1_33to32:writedata
	signal irq_mapper_receiver0_irq                                                  : std_logic;                     -- epcs_flash_controller:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                  : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                               : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                            : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                        : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, epcs_flash_controller:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                             : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in1
	signal reset_n_reset_n_ports_inv                                                 : std_logic;                     -- reset_n_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv              : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv             : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_0_epcs_flash_controller_epcs_control_port_read:inv -> epcs_flash_controller:read_n
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_0_epcs_flash_controller_epcs_control_port_write:inv -> epcs_flash_controller:write_n
	signal mm_interconnect_0_po_led_s1_write_ports_inv                               : std_logic;                     -- mm_interconnect_0_po_led_s1_write:inv -> po_led:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                                 : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                                : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_pio_gpio2_s1_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_pio_gpio2_s1_write:inv -> pio_gpio2:write_n
	signal mm_interconnect_0_pio_gpio0_31to0_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_pio_gpio0_31to0_s1_write:inv -> pio_gpio0_31to0:write_n
	signal mm_interconnect_0_pio_gpio1_31to0_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_pio_gpio1_31to0_s1_write:inv -> pio_gpio1_31to0:write_n
	signal mm_interconnect_0_pio_gpio0_33to32_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_pio_gpio0_33to32_s1_write:inv -> pio_gpio0_33to32:write_n
	signal mm_interconnect_0_pio_gpio1_33to32_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_pio_gpio1_33to32_s1_write:inv -> pio_gpio1_33to32:write_n
	signal rst_controller_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, epcs_flash_controller:reset_n, jtag_uart:rst_n, pi_gpio0:reset_n, pi_gpio1:reset_n, pi_gpio2:reset_n, pi_key:reset_n, pi_sw:reset_n, pio_gpio0_31to0:reset_n, pio_gpio0_33to32:reset_n, pio_gpio1_31to0:reset_n, pio_gpio1_33to32:reset_n, pio_gpio2:reset_n, po_led:reset_n, sdram:reset_n, sysid:reset_n]

begin

	cpu : component crypto_wallet_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	epcs_flash_controller : component crypto_wallet_epcs_flash_controller
		port map (
			clk        => clk_clk,                                                                   --               clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                                  --             reset.reset_n
			reset_req  => rst_controller_reset_out_reset_req,                                        --                  .reset_req
			address    => mm_interconnect_0_epcs_flash_controller_epcs_control_port_address,         -- epcs_control_port.address
			chipselect => mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect,      --                  .chipselect
			read_n     => mm_interconnect_0_epcs_flash_controller_epcs_control_port_read_ports_inv,  --                  .read_n
			readdata   => mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata,        --                  .readdata
			write_n    => mm_interconnect_0_epcs_flash_controller_epcs_control_port_write_ports_inv, --                  .write_n
			writedata  => mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata,       --                  .writedata
			irq        => irq_mapper_receiver0_irq,                                                  --               irq.irq
			dclk       => epcs_flash_controller_dclk,                                                --          external.export
			sce        => epcs_flash_controller_sce,                                                 --                  .export
			sdo        => epcs_flash_controller_sdo,                                                 --                  .export
			data0      => epcs_flash_controller_data0                                                --                  .export
		);

	jtag_uart : component crypto_wallet_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	onchip_memory2 : component crypto_wallet_onchip_memory2
		port map (
			clk        => clk_clk,                                        --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,             --       .reset_req
			freeze     => '0'                                             -- (terminated)
		);

	pi_gpio0 : component crypto_wallet_pi_gpio0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pi_gpio0_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_pi_gpio0_s1_readdata,   --                    .readdata
			in_port  => pi_gpio0_external_connection_export       -- external_connection.export
		);

	pi_gpio1 : component crypto_wallet_pi_gpio0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pi_gpio1_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_pi_gpio1_s1_readdata,   --                    .readdata
			in_port  => pi_gpio1_external_connection_export       -- external_connection.export
		);

	pi_gpio2 : component crypto_wallet_pi_gpio2
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pi_gpio2_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_pi_gpio2_s1_readdata,   --                    .readdata
			in_port  => pi_gpio2_external_connection_export       -- external_connection.export
		);

	pi_key : component crypto_wallet_pi_gpio0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pi_key_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_pi_key_s1_readdata,     --                    .readdata
			in_port  => pi_key_external_connection_export         -- external_connection.export
		);

	pi_sw : component crypto_wallet_pi_sw
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pi_sw_s1_address,       --                  s1.address
			readdata => mm_interconnect_0_pi_sw_s1_readdata,      --                    .readdata
			in_port  => pi_sw_external_connection_export          -- external_connection.export
		);

	pio_gpio0_31to0 : component crypto_wallet_pio_gpio0_31to0
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_pio_gpio0_31to0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_gpio0_31to0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_gpio0_31to0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_gpio0_31to0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_gpio0_31to0_s1_readdata,        --                    .readdata
			bidir_port => pio_gpio0_external_connection_export                  -- external_connection.export
		);

	pio_gpio0_33to32 : component crypto_wallet_pio_gpio0_33to32
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_pio_gpio0_33to32_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_gpio0_33to32_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_gpio0_33to32_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_gpio0_33to32_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_gpio0_33to32_s1_readdata,        --                    .readdata
			bidir_port => pio_gpio0_33to32_external_connection_export            -- external_connection.export
		);

	pio_gpio1_31to0 : component crypto_wallet_pio_gpio0_31to0
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_pio_gpio1_31to0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_gpio1_31to0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_gpio1_31to0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_gpio1_31to0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_gpio1_31to0_s1_readdata,        --                    .readdata
			bidir_port => pio_gpio1_external_connection_export                  -- external_connection.export
		);

	pio_gpio1_33to32 : component crypto_wallet_pio_gpio0_33to32
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_pio_gpio1_33to32_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_gpio1_33to32_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_gpio1_33to32_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_gpio1_33to32_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_gpio1_33to32_s1_readdata,        --                    .readdata
			bidir_port => pio_gpio1_33to32_external_connection_export            -- external_connection.export
		);

	pio_gpio2 : component crypto_wallet_pio_gpio2
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_pio_gpio2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_gpio2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_gpio2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_gpio2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_gpio2_s1_readdata,        --                    .readdata
			bidir_port => pio_gpio2_external_connection_export            -- external_connection.export
		);

	po_led : component crypto_wallet_po_led
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_po_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_po_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_po_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_po_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_po_led_s1_readdata,        --                    .readdata
			out_port   => po_led_external_connection_export            -- external_connection.export
		);

	sdram : component crypto_wallet_sdram
		port map (
			clk            => clk_clk,                                         --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	sysid : component crypto_wallet_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component crypto_wallet_mm_interconnect_0
		port map (
			clk_50_clk_clk                                     => clk_clk,                                                              --                              clk_50_clk.clk
			cpu_reset_reset_bridge_in_reset_reset              => rst_controller_reset_out_reset,                                       --         cpu_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                            => cpu_data_master_address,                                              --                         cpu_data_master.address
			cpu_data_master_waitrequest                        => cpu_data_master_waitrequest,                                          --                                        .waitrequest
			cpu_data_master_byteenable                         => cpu_data_master_byteenable,                                           --                                        .byteenable
			cpu_data_master_read                               => cpu_data_master_read,                                                 --                                        .read
			cpu_data_master_readdata                           => cpu_data_master_readdata,                                             --                                        .readdata
			cpu_data_master_write                              => cpu_data_master_write,                                                --                                        .write
			cpu_data_master_writedata                          => cpu_data_master_writedata,                                            --                                        .writedata
			cpu_data_master_debugaccess                        => cpu_data_master_debugaccess,                                          --                                        .debugaccess
			cpu_instruction_master_address                     => cpu_instruction_master_address,                                       --                  cpu_instruction_master.address
			cpu_instruction_master_waitrequest                 => cpu_instruction_master_waitrequest,                                   --                                        .waitrequest
			cpu_instruction_master_read                        => cpu_instruction_master_read,                                          --                                        .read
			cpu_instruction_master_readdata                    => cpu_instruction_master_readdata,                                      --                                        .readdata
			cpu_debug_mem_slave_address                        => mm_interconnect_0_cpu_debug_mem_slave_address,                        --                     cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                          => mm_interconnect_0_cpu_debug_mem_slave_write,                          --                                        .write
			cpu_debug_mem_slave_read                           => mm_interconnect_0_cpu_debug_mem_slave_read,                           --                                        .read
			cpu_debug_mem_slave_readdata                       => mm_interconnect_0_cpu_debug_mem_slave_readdata,                       --                                        .readdata
			cpu_debug_mem_slave_writedata                      => mm_interconnect_0_cpu_debug_mem_slave_writedata,                      --                                        .writedata
			cpu_debug_mem_slave_byteenable                     => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                     --                                        .byteenable
			cpu_debug_mem_slave_waitrequest                    => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                    --                                        .waitrequest
			cpu_debug_mem_slave_debugaccess                    => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                    --                                        .debugaccess
			epcs_flash_controller_epcs_control_port_address    => mm_interconnect_0_epcs_flash_controller_epcs_control_port_address,    -- epcs_flash_controller_epcs_control_port.address
			epcs_flash_controller_epcs_control_port_write      => mm_interconnect_0_epcs_flash_controller_epcs_control_port_write,      --                                        .write
			epcs_flash_controller_epcs_control_port_read       => mm_interconnect_0_epcs_flash_controller_epcs_control_port_read,       --                                        .read
			epcs_flash_controller_epcs_control_port_readdata   => mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata,   --                                        .readdata
			epcs_flash_controller_epcs_control_port_writedata  => mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata,  --                                        .writedata
			epcs_flash_controller_epcs_control_port_chipselect => mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect, --                                        .chipselect
			jtag_uart_avalon_jtag_slave_address                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,                --             jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                  --                                        .write
			jtag_uart_avalon_jtag_slave_read                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                   --                                        .read
			jtag_uart_avalon_jtag_slave_readdata               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,               --                                        .readdata
			jtag_uart_avalon_jtag_slave_writedata              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,              --                                        .writedata
			jtag_uart_avalon_jtag_slave_waitrequest            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,            --                                        .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,             --                                        .chipselect
			onchip_memory2_s1_address                          => mm_interconnect_0_onchip_memory2_s1_address,                          --                       onchip_memory2_s1.address
			onchip_memory2_s1_write                            => mm_interconnect_0_onchip_memory2_s1_write,                            --                                        .write
			onchip_memory2_s1_readdata                         => mm_interconnect_0_onchip_memory2_s1_readdata,                         --                                        .readdata
			onchip_memory2_s1_writedata                        => mm_interconnect_0_onchip_memory2_s1_writedata,                        --                                        .writedata
			onchip_memory2_s1_byteenable                       => mm_interconnect_0_onchip_memory2_s1_byteenable,                       --                                        .byteenable
			onchip_memory2_s1_chipselect                       => mm_interconnect_0_onchip_memory2_s1_chipselect,                       --                                        .chipselect
			onchip_memory2_s1_clken                            => mm_interconnect_0_onchip_memory2_s1_clken,                            --                                        .clken
			pi_gpio0_s1_address                                => mm_interconnect_0_pi_gpio0_s1_address,                                --                             pi_gpio0_s1.address
			pi_gpio0_s1_readdata                               => mm_interconnect_0_pi_gpio0_s1_readdata,                               --                                        .readdata
			pi_gpio1_s1_address                                => mm_interconnect_0_pi_gpio1_s1_address,                                --                             pi_gpio1_s1.address
			pi_gpio1_s1_readdata                               => mm_interconnect_0_pi_gpio1_s1_readdata,                               --                                        .readdata
			pi_gpio2_s1_address                                => mm_interconnect_0_pi_gpio2_s1_address,                                --                             pi_gpio2_s1.address
			pi_gpio2_s1_readdata                               => mm_interconnect_0_pi_gpio2_s1_readdata,                               --                                        .readdata
			pi_key_s1_address                                  => mm_interconnect_0_pi_key_s1_address,                                  --                               pi_key_s1.address
			pi_key_s1_readdata                                 => mm_interconnect_0_pi_key_s1_readdata,                                 --                                        .readdata
			pi_sw_s1_address                                   => mm_interconnect_0_pi_sw_s1_address,                                   --                                pi_sw_s1.address
			pi_sw_s1_readdata                                  => mm_interconnect_0_pi_sw_s1_readdata,                                  --                                        .readdata
			pio_gpio0_31to0_s1_address                         => mm_interconnect_0_pio_gpio0_31to0_s1_address,                         --                      pio_gpio0_31to0_s1.address
			pio_gpio0_31to0_s1_write                           => mm_interconnect_0_pio_gpio0_31to0_s1_write,                           --                                        .write
			pio_gpio0_31to0_s1_readdata                        => mm_interconnect_0_pio_gpio0_31to0_s1_readdata,                        --                                        .readdata
			pio_gpio0_31to0_s1_writedata                       => mm_interconnect_0_pio_gpio0_31to0_s1_writedata,                       --                                        .writedata
			pio_gpio0_31to0_s1_chipselect                      => mm_interconnect_0_pio_gpio0_31to0_s1_chipselect,                      --                                        .chipselect
			pio_gpio0_33to32_s1_address                        => mm_interconnect_0_pio_gpio0_33to32_s1_address,                        --                     pio_gpio0_33to32_s1.address
			pio_gpio0_33to32_s1_write                          => mm_interconnect_0_pio_gpio0_33to32_s1_write,                          --                                        .write
			pio_gpio0_33to32_s1_readdata                       => mm_interconnect_0_pio_gpio0_33to32_s1_readdata,                       --                                        .readdata
			pio_gpio0_33to32_s1_writedata                      => mm_interconnect_0_pio_gpio0_33to32_s1_writedata,                      --                                        .writedata
			pio_gpio0_33to32_s1_chipselect                     => mm_interconnect_0_pio_gpio0_33to32_s1_chipselect,                     --                                        .chipselect
			pio_gpio1_31to0_s1_address                         => mm_interconnect_0_pio_gpio1_31to0_s1_address,                         --                      pio_gpio1_31to0_s1.address
			pio_gpio1_31to0_s1_write                           => mm_interconnect_0_pio_gpio1_31to0_s1_write,                           --                                        .write
			pio_gpio1_31to0_s1_readdata                        => mm_interconnect_0_pio_gpio1_31to0_s1_readdata,                        --                                        .readdata
			pio_gpio1_31to0_s1_writedata                       => mm_interconnect_0_pio_gpio1_31to0_s1_writedata,                       --                                        .writedata
			pio_gpio1_31to0_s1_chipselect                      => mm_interconnect_0_pio_gpio1_31to0_s1_chipselect,                      --                                        .chipselect
			pio_gpio1_33to32_s1_address                        => mm_interconnect_0_pio_gpio1_33to32_s1_address,                        --                     pio_gpio1_33to32_s1.address
			pio_gpio1_33to32_s1_write                          => mm_interconnect_0_pio_gpio1_33to32_s1_write,                          --                                        .write
			pio_gpio1_33to32_s1_readdata                       => mm_interconnect_0_pio_gpio1_33to32_s1_readdata,                       --                                        .readdata
			pio_gpio1_33to32_s1_writedata                      => mm_interconnect_0_pio_gpio1_33to32_s1_writedata,                      --                                        .writedata
			pio_gpio1_33to32_s1_chipselect                     => mm_interconnect_0_pio_gpio1_33to32_s1_chipselect,                     --                                        .chipselect
			pio_gpio2_s1_address                               => mm_interconnect_0_pio_gpio2_s1_address,                               --                            pio_gpio2_s1.address
			pio_gpio2_s1_write                                 => mm_interconnect_0_pio_gpio2_s1_write,                                 --                                        .write
			pio_gpio2_s1_readdata                              => mm_interconnect_0_pio_gpio2_s1_readdata,                              --                                        .readdata
			pio_gpio2_s1_writedata                             => mm_interconnect_0_pio_gpio2_s1_writedata,                             --                                        .writedata
			pio_gpio2_s1_chipselect                            => mm_interconnect_0_pio_gpio2_s1_chipselect,                            --                                        .chipselect
			po_led_s1_address                                  => mm_interconnect_0_po_led_s1_address,                                  --                               po_led_s1.address
			po_led_s1_write                                    => mm_interconnect_0_po_led_s1_write,                                    --                                        .write
			po_led_s1_readdata                                 => mm_interconnect_0_po_led_s1_readdata,                                 --                                        .readdata
			po_led_s1_writedata                                => mm_interconnect_0_po_led_s1_writedata,                                --                                        .writedata
			po_led_s1_chipselect                               => mm_interconnect_0_po_led_s1_chipselect,                               --                                        .chipselect
			sdram_s1_address                                   => mm_interconnect_0_sdram_s1_address,                                   --                                sdram_s1.address
			sdram_s1_write                                     => mm_interconnect_0_sdram_s1_write,                                     --                                        .write
			sdram_s1_read                                      => mm_interconnect_0_sdram_s1_read,                                      --                                        .read
			sdram_s1_readdata                                  => mm_interconnect_0_sdram_s1_readdata,                                  --                                        .readdata
			sdram_s1_writedata                                 => mm_interconnect_0_sdram_s1_writedata,                                 --                                        .writedata
			sdram_s1_byteenable                                => mm_interconnect_0_sdram_s1_byteenable,                                --                                        .byteenable
			sdram_s1_readdatavalid                             => mm_interconnect_0_sdram_s1_readdatavalid,                             --                                        .readdatavalid
			sdram_s1_waitrequest                               => mm_interconnect_0_sdram_s1_waitrequest,                               --                                        .waitrequest
			sdram_s1_chipselect                                => mm_interconnect_0_sdram_s1_chipselect,                                --                                        .chipselect
			sysid_control_slave_address                        => mm_interconnect_0_sysid_control_slave_address,                        --                     sysid_control_slave.address
			sysid_control_slave_readdata                       => mm_interconnect_0_sysid_control_slave_readdata                        --                                        .readdata
		);

	irq_mapper : component crypto_wallet_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_n_reset_n_ports_inv,          -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_n_reset_n_ports_inv <= not reset_n_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_epcs_flash_controller_epcs_control_port_read_ports_inv <= not mm_interconnect_0_epcs_flash_controller_epcs_control_port_read;

	mm_interconnect_0_epcs_flash_controller_epcs_control_port_write_ports_inv <= not mm_interconnect_0_epcs_flash_controller_epcs_control_port_write;

	mm_interconnect_0_po_led_s1_write_ports_inv <= not mm_interconnect_0_po_led_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_pio_gpio2_s1_write_ports_inv <= not mm_interconnect_0_pio_gpio2_s1_write;

	mm_interconnect_0_pio_gpio0_31to0_s1_write_ports_inv <= not mm_interconnect_0_pio_gpio0_31to0_s1_write;

	mm_interconnect_0_pio_gpio1_31to0_s1_write_ports_inv <= not mm_interconnect_0_pio_gpio1_31to0_s1_write;

	mm_interconnect_0_pio_gpio0_33to32_s1_write_ports_inv <= not mm_interconnect_0_pio_gpio0_33to32_s1_write;

	mm_interconnect_0_pio_gpio1_33to32_s1_write_ports_inv <= not mm_interconnect_0_pio_gpio1_33to32_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of crypto_wallet
