// crypto_wallet2_nios.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module crypto_wallet2_nios (
		input  wire        clk_clk,                                      //                                   clk.clk
		output wire        epcs_flash_controller_external_dclk,          //        epcs_flash_controller_external.dclk
		output wire        epcs_flash_controller_external_sce,           //                                      .sce
		output wire        epcs_flash_controller_external_sdo,           //                                      .sdo
		input  wire        epcs_flash_controller_external_data0,         //                                      .data0
		input  wire [7:0]  pi_random_external_connection_export,         //         pi_random_external_connection.export
		output wire [7:0]  po_led_external_connection_export,            //            po_led_external_connection.export
		output wire [31:0] po_random_seed_external_connection_export,    //    po_random_seed_external_connection.export
		output wire [7:0]  po_system_control_external_connection_export, // po_system_control_external_connection.export
		input  wire        reset_reset_n,                                //                                 reset.reset_n
		output wire [12:0] sdram_wire_addr,                              //                            sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                //                                      .ba
		output wire        sdram_wire_cas_n,                             //                                      .cas_n
		output wire        sdram_wire_cke,                               //                                      .cke
		output wire        sdram_wire_cs_n,                              //                                      .cs_n
		inout  wire [15:0] sdram_wire_dq,                                //                                      .dq
		output wire [1:0]  sdram_wire_dqm,                               //                                      .dqm
		output wire        sdram_wire_ras_n,                             //                                      .ras_n
		output wire        sdram_wire_we_n,                              //                                      .we_n
		input  wire        uart_external_connection_rxd,                 //              uart_external_connection.rxd
		output wire        uart_external_connection_txd                  //                                      .txd
	);

	wire  [31:0] cpu_data_master_readdata;                                             // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                          // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                          // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [25:0] cpu_data_master_address;                                              // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                           // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                 // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                                // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                            // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                      // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                   // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [25:0] cpu_instruction_master_address;                                       // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                          // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;               // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;            // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                       // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                        // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                       // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                    // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                    // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                        // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                           // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                     // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                          // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                      // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_controller_epcs_control_port_chipselect -> epcs_flash_controller:chipselect
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata;   // epcs_flash_controller:readdata -> mm_interconnect_0:epcs_flash_controller_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_controller_epcs_control_port_address -> epcs_flash_controller:address
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_controller_epcs_control_port_read -> epcs_flash_controller:read_n
	wire         mm_interconnect_0_epcs_flash_controller_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_controller_epcs_control_port_write -> epcs_flash_controller:write_n
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_controller_epcs_control_port_writedata -> epcs_flash_controller:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                       // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                         // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_s1_address;                          // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                       // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                            // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                        // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                            // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_po_led_s1_chipselect;                               // mm_interconnect_0:po_led_s1_chipselect -> po_led:chipselect
	wire  [31:0] mm_interconnect_0_po_led_s1_readdata;                                 // po_led:readdata -> mm_interconnect_0:po_led_s1_readdata
	wire   [1:0] mm_interconnect_0_po_led_s1_address;                                  // mm_interconnect_0:po_led_s1_address -> po_led:address
	wire         mm_interconnect_0_po_led_s1_write;                                    // mm_interconnect_0:po_led_s1_write -> po_led:write_n
	wire  [31:0] mm_interconnect_0_po_led_s1_writedata;                                // mm_interconnect_0:po_led_s1_writedata -> po_led:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                  // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                               // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                   // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                      // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                             // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                     // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                 // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_uart_s1_chipselect;                                 // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                                   // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                                    // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                                       // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                              // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                                      // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                                  // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire  [31:0] mm_interconnect_0_pi_random_value_s1_readdata;                        // pi_random_value:readdata -> mm_interconnect_0:pi_random_value_s1_readdata
	wire   [1:0] mm_interconnect_0_pi_random_value_s1_address;                         // mm_interconnect_0:pi_random_value_s1_address -> pi_random_value:address
	wire         mm_interconnect_0_po_system_control_s1_chipselect;                    // mm_interconnect_0:po_system_control_s1_chipselect -> po_system_control:chipselect
	wire  [31:0] mm_interconnect_0_po_system_control_s1_readdata;                      // po_system_control:readdata -> mm_interconnect_0:po_system_control_s1_readdata
	wire   [1:0] mm_interconnect_0_po_system_control_s1_address;                       // mm_interconnect_0:po_system_control_s1_address -> po_system_control:address
	wire         mm_interconnect_0_po_system_control_s1_write;                         // mm_interconnect_0:po_system_control_s1_write -> po_system_control:write_n
	wire  [31:0] mm_interconnect_0_po_system_control_s1_writedata;                     // mm_interconnect_0:po_system_control_s1_writedata -> po_system_control:writedata
	wire         mm_interconnect_0_po_random_seed_s1_chipselect;                       // mm_interconnect_0:po_random_seed_s1_chipselect -> po_random_seed:chipselect
	wire  [31:0] mm_interconnect_0_po_random_seed_s1_readdata;                         // po_random_seed:readdata -> mm_interconnect_0:po_random_seed_s1_readdata
	wire   [1:0] mm_interconnect_0_po_random_seed_s1_address;                          // mm_interconnect_0:po_random_seed_s1_address -> po_random_seed:address
	wire         mm_interconnect_0_po_random_seed_s1_write;                            // mm_interconnect_0:po_random_seed_s1_write -> po_random_seed:write_n
	wire  [31:0] mm_interconnect_0_po_random_seed_s1_writedata;                        // mm_interconnect_0:po_random_seed_s1_writedata -> po_random_seed:writedata
	wire         irq_mapper_receiver0_irq;                                             // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                             // epcs_flash_controller:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                             // uart:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                                          // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_reset_out_reset_req;                                   // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                        // cpu:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [epcs_flash_controller:reset_n, jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, pi_random_value:reset_n, po_led:reset_n, po_random_seed:reset_n, po_system_control:reset_n, rst_translator_001:in_reset, sdram:reset_n, sysid:reset_n, uart:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                               // rst_controller_001:reset_req -> [epcs_flash_controller:reset_req, onchip_memory2:reset_req, rst_translator_001:reset_req_in]

	crypto_wallet2_nios_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	crypto_wallet2_nios_epcs_flash_controller epcs_flash_controller (
		.clk        (clk_clk),                                                              //               clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                                  //             reset.reset_n
		.reset_req  (rst_controller_001_reset_out_reset_req),                               //                  .reset_req
		.address    (mm_interconnect_0_epcs_flash_controller_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_flash_controller_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_flash_controller_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver1_irq),                                             //               irq.irq
		.dclk       (epcs_flash_controller_external_dclk),                                  //          external.export
		.sce        (epcs_flash_controller_external_sce),                                   //                  .export
		.sdo        (epcs_flash_controller_external_sdo),                                   //                  .export
		.data0      (epcs_flash_controller_external_data0)                                  //                  .export
	);

	crypto_wallet2_nios_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	crypto_wallet2_nios_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	crypto_wallet2_nios_pi_random_value pi_random_value (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_pi_random_value_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pi_random_value_s1_readdata), //                    .readdata
		.in_port  (pi_random_external_connection_export)           // external_connection.export
	);

	crypto_wallet2_nios_po_led po_led (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_po_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_led_s1_readdata),   //                    .readdata
		.out_port   (po_led_external_connection_export)       // external_connection.export
	);

	crypto_wallet2_nios_po_random_seed po_random_seed (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_po_random_seed_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_random_seed_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_random_seed_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_random_seed_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_random_seed_s1_readdata),   //                    .readdata
		.out_port   (po_random_seed_external_connection_export)       // external_connection.export
	);

	crypto_wallet2_nios_po_led po_system_control (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_po_system_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_po_system_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_po_system_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_po_system_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_po_system_control_s1_readdata),   //                    .readdata
		.out_port   (po_system_control_external_connection_export)       // external_connection.export
	);

	crypto_wallet2_nios_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	crypto_wallet2_nios_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	crypto_wallet2_nios_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_external_connection_rxd),            // external_connection.export
		.txd           (uart_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	crypto_wallet2_nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                     (clk_clk),                                                              //                              clk_50_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                                       //         cpu_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                                   //   jtag_uart_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                            (cpu_data_master_address),                                              //                         cpu_data_master.address
		.cpu_data_master_waitrequest                        (cpu_data_master_waitrequest),                                          //                                        .waitrequest
		.cpu_data_master_byteenable                         (cpu_data_master_byteenable),                                           //                                        .byteenable
		.cpu_data_master_read                               (cpu_data_master_read),                                                 //                                        .read
		.cpu_data_master_readdata                           (cpu_data_master_readdata),                                             //                                        .readdata
		.cpu_data_master_write                              (cpu_data_master_write),                                                //                                        .write
		.cpu_data_master_writedata                          (cpu_data_master_writedata),                                            //                                        .writedata
		.cpu_data_master_debugaccess                        (cpu_data_master_debugaccess),                                          //                                        .debugaccess
		.cpu_instruction_master_address                     (cpu_instruction_master_address),                                       //                  cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                 (cpu_instruction_master_waitrequest),                                   //                                        .waitrequest
		.cpu_instruction_master_read                        (cpu_instruction_master_read),                                          //                                        .read
		.cpu_instruction_master_readdata                    (cpu_instruction_master_readdata),                                      //                                        .readdata
		.cpu_debug_mem_slave_address                        (mm_interconnect_0_cpu_debug_mem_slave_address),                        //                     cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                          (mm_interconnect_0_cpu_debug_mem_slave_write),                          //                                        .write
		.cpu_debug_mem_slave_read                           (mm_interconnect_0_cpu_debug_mem_slave_read),                           //                                        .read
		.cpu_debug_mem_slave_readdata                       (mm_interconnect_0_cpu_debug_mem_slave_readdata),                       //                                        .readdata
		.cpu_debug_mem_slave_writedata                      (mm_interconnect_0_cpu_debug_mem_slave_writedata),                      //                                        .writedata
		.cpu_debug_mem_slave_byteenable                     (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                     //                                        .byteenable
		.cpu_debug_mem_slave_waitrequest                    (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                    //                                        .waitrequest
		.cpu_debug_mem_slave_debugaccess                    (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                    //                                        .debugaccess
		.epcs_flash_controller_epcs_control_port_address    (mm_interconnect_0_epcs_flash_controller_epcs_control_port_address),    // epcs_flash_controller_epcs_control_port.address
		.epcs_flash_controller_epcs_control_port_write      (mm_interconnect_0_epcs_flash_controller_epcs_control_port_write),      //                                        .write
		.epcs_flash_controller_epcs_control_port_read       (mm_interconnect_0_epcs_flash_controller_epcs_control_port_read),       //                                        .read
		.epcs_flash_controller_epcs_control_port_readdata   (mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata),   //                                        .readdata
		.epcs_flash_controller_epcs_control_port_writedata  (mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata),  //                                        .writedata
		.epcs_flash_controller_epcs_control_port_chipselect (mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect), //                                        .chipselect
		.jtag_uart_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                //             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                  //                                        .write
		.jtag_uart_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                   //                                        .read
		.jtag_uart_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),               //                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),              //                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),            //                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),             //                                        .chipselect
		.onchip_memory2_s1_address                          (mm_interconnect_0_onchip_memory2_s1_address),                          //                       onchip_memory2_s1.address
		.onchip_memory2_s1_write                            (mm_interconnect_0_onchip_memory2_s1_write),                            //                                        .write
		.onchip_memory2_s1_readdata                         (mm_interconnect_0_onchip_memory2_s1_readdata),                         //                                        .readdata
		.onchip_memory2_s1_writedata                        (mm_interconnect_0_onchip_memory2_s1_writedata),                        //                                        .writedata
		.onchip_memory2_s1_byteenable                       (mm_interconnect_0_onchip_memory2_s1_byteenable),                       //                                        .byteenable
		.onchip_memory2_s1_chipselect                       (mm_interconnect_0_onchip_memory2_s1_chipselect),                       //                                        .chipselect
		.onchip_memory2_s1_clken                            (mm_interconnect_0_onchip_memory2_s1_clken),                            //                                        .clken
		.pi_random_value_s1_address                         (mm_interconnect_0_pi_random_value_s1_address),                         //                      pi_random_value_s1.address
		.pi_random_value_s1_readdata                        (mm_interconnect_0_pi_random_value_s1_readdata),                        //                                        .readdata
		.po_led_s1_address                                  (mm_interconnect_0_po_led_s1_address),                                  //                               po_led_s1.address
		.po_led_s1_write                                    (mm_interconnect_0_po_led_s1_write),                                    //                                        .write
		.po_led_s1_readdata                                 (mm_interconnect_0_po_led_s1_readdata),                                 //                                        .readdata
		.po_led_s1_writedata                                (mm_interconnect_0_po_led_s1_writedata),                                //                                        .writedata
		.po_led_s1_chipselect                               (mm_interconnect_0_po_led_s1_chipselect),                               //                                        .chipselect
		.po_random_seed_s1_address                          (mm_interconnect_0_po_random_seed_s1_address),                          //                       po_random_seed_s1.address
		.po_random_seed_s1_write                            (mm_interconnect_0_po_random_seed_s1_write),                            //                                        .write
		.po_random_seed_s1_readdata                         (mm_interconnect_0_po_random_seed_s1_readdata),                         //                                        .readdata
		.po_random_seed_s1_writedata                        (mm_interconnect_0_po_random_seed_s1_writedata),                        //                                        .writedata
		.po_random_seed_s1_chipselect                       (mm_interconnect_0_po_random_seed_s1_chipselect),                       //                                        .chipselect
		.po_system_control_s1_address                       (mm_interconnect_0_po_system_control_s1_address),                       //                    po_system_control_s1.address
		.po_system_control_s1_write                         (mm_interconnect_0_po_system_control_s1_write),                         //                                        .write
		.po_system_control_s1_readdata                      (mm_interconnect_0_po_system_control_s1_readdata),                      //                                        .readdata
		.po_system_control_s1_writedata                     (mm_interconnect_0_po_system_control_s1_writedata),                     //                                        .writedata
		.po_system_control_s1_chipselect                    (mm_interconnect_0_po_system_control_s1_chipselect),                    //                                        .chipselect
		.sdram_s1_address                                   (mm_interconnect_0_sdram_s1_address),                                   //                                sdram_s1.address
		.sdram_s1_write                                     (mm_interconnect_0_sdram_s1_write),                                     //                                        .write
		.sdram_s1_read                                      (mm_interconnect_0_sdram_s1_read),                                      //                                        .read
		.sdram_s1_readdata                                  (mm_interconnect_0_sdram_s1_readdata),                                  //                                        .readdata
		.sdram_s1_writedata                                 (mm_interconnect_0_sdram_s1_writedata),                                 //                                        .writedata
		.sdram_s1_byteenable                                (mm_interconnect_0_sdram_s1_byteenable),                                //                                        .byteenable
		.sdram_s1_readdatavalid                             (mm_interconnect_0_sdram_s1_readdatavalid),                             //                                        .readdatavalid
		.sdram_s1_waitrequest                               (mm_interconnect_0_sdram_s1_waitrequest),                               //                                        .waitrequest
		.sdram_s1_chipselect                                (mm_interconnect_0_sdram_s1_chipselect),                                //                                        .chipselect
		.sysid_control_slave_address                        (mm_interconnect_0_sysid_control_slave_address),                        //                     sysid_control_slave.address
		.sysid_control_slave_readdata                       (mm_interconnect_0_sysid_control_slave_readdata),                       //                                        .readdata
		.uart_s1_address                                    (mm_interconnect_0_uart_s1_address),                                    //                                 uart_s1.address
		.uart_s1_write                                      (mm_interconnect_0_uart_s1_write),                                      //                                        .write
		.uart_s1_read                                       (mm_interconnect_0_uart_s1_read),                                       //                                        .read
		.uart_s1_readdata                                   (mm_interconnect_0_uart_s1_readdata),                                   //                                        .readdata
		.uart_s1_writedata                                  (mm_interconnect_0_uart_s1_writedata),                                  //                                        .writedata
		.uart_s1_begintransfer                              (mm_interconnect_0_uart_s1_begintransfer),                              //                                        .begintransfer
		.uart_s1_chipselect                                 (mm_interconnect_0_uart_s1_chipselect)                                  //                                        .chipselect
	);

	crypto_wallet2_nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
