-- crypto_wallet.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity crypto_wallet is
	port (
		buttons_pi_export : in    std_logic_vector(1 downto 0)  := (others => '0'); -- buttons_pi.export
		clk_clk           : in    std_logic                     := '0';             --        clk.clk
		epcs_dclk         : out   std_logic;                                        --       epcs.dclk
		epcs_sce          : out   std_logic;                                        --           .sce
		epcs_sdo          : out   std_logic;                                        --           .sdo
		epcs_data0        : in    std_logic                     := '0';             --           .data0
		led_po_export     : out   std_logic_vector(7 downto 0);                     --     led_po.export
		reset_reset_n     : in    std_logic                     := '0';             --      reset.reset_n
		sdram_addr        : out   std_logic_vector(12 downto 0);                    --      sdram.addr
		sdram_ba          : out   std_logic_vector(1 downto 0);                     --           .ba
		sdram_cas_n       : out   std_logic;                                        --           .cas_n
		sdram_cke         : out   std_logic;                                        --           .cke
		sdram_cs_n        : out   std_logic;                                        --           .cs_n
		sdram_dq          : inout std_logic_vector(15 downto 0) := (others => '0'); --           .dq
		sdram_dqm         : out   std_logic_vector(1 downto 0);                     --           .dqm
		sdram_ras_n       : out   std_logic;                                        --           .ras_n
		sdram_we_n        : out   std_logic;                                        --           .we_n
		switch_pi_export  : in    std_logic_vector(3 downto 0)  := (others => '0'); --  switch_pi.export
		uart_0_rxd        : in    std_logic                     := '0';             --     uart_0.rxd
		uart_0_txd        : out   std_logic                                         --           .txd
	);
end entity crypto_wallet;

architecture rtl of crypto_wallet is
	component crypto_wallet_buttons_pi is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			KEY        : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component crypto_wallet_buttons_pi;

	component crypto_wallet_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component crypto_wallet_cpu;

	component crypto_wallet_epcs_flash_controller is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read_n     : in  std_logic                     := 'X';             -- read_n
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq        : out std_logic;                                        -- irq
			dclk       : out std_logic;                                        -- export
			sce        : out std_logic;                                        -- export
			sdo        : out std_logic;                                        -- export
			data0      : in  std_logic                     := 'X'              -- export
		);
	end component crypto_wallet_epcs_flash_controller;

	component crypto_wallet_led_po is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			LEDG       : out std_logic_vector(7 downto 0)                      -- export
		);
	end component crypto_wallet_led_po;

	component crypto_wallet_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component crypto_wallet_sdram;

	component crypto_wallet_switch_pi is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			DIP        : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component crypto_wallet_switch_pi;

	component crypto_wallet_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component crypto_wallet_sysid;

	component crypto_wallet_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component crypto_wallet_uart_0;

	component crypto_wallet_mm_interconnect_0 is
		port (
			clk_sys_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                            : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                        : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                               : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                              : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                        : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                 : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                        : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			buttons_pi_avalon_parallel_port_slave_address      : out std_logic_vector(1 downto 0);                     -- address
			buttons_pi_avalon_parallel_port_slave_write        : out std_logic;                                        -- write
			buttons_pi_avalon_parallel_port_slave_read         : out std_logic;                                        -- read
			buttons_pi_avalon_parallel_port_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			buttons_pi_avalon_parallel_port_slave_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			buttons_pi_avalon_parallel_port_slave_byteenable   : out std_logic_vector(3 downto 0);                     -- byteenable
			buttons_pi_avalon_parallel_port_slave_chipselect   : out std_logic;                                        -- chipselect
			cpu_debug_mem_slave_address                        : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                          : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                           : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                    : out std_logic;                                        -- debugaccess
			epcs_flash_controller_epcs_control_port_address    : out std_logic_vector(8 downto 0);                     -- address
			epcs_flash_controller_epcs_control_port_write      : out std_logic;                                        -- write
			epcs_flash_controller_epcs_control_port_read       : out std_logic;                                        -- read
			epcs_flash_controller_epcs_control_port_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			epcs_flash_controller_epcs_control_port_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			epcs_flash_controller_epcs_control_port_chipselect : out std_logic;                                        -- chipselect
			led_po_avalon_parallel_port_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			led_po_avalon_parallel_port_slave_write            : out std_logic;                                        -- write
			led_po_avalon_parallel_port_slave_read             : out std_logic;                                        -- read
			led_po_avalon_parallel_port_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_po_avalon_parallel_port_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			led_po_avalon_parallel_port_slave_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			led_po_avalon_parallel_port_slave_chipselect       : out std_logic;                                        -- chipselect
			sdram_s1_address                                   : out std_logic_vector(23 downto 0);                    -- address
			sdram_s1_write                                     : out std_logic;                                        -- write
			sdram_s1_read                                      : out std_logic;                                        -- read
			sdram_s1_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                             : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                : out std_logic;                                        -- chipselect
			switch_pi_avalon_parallel_port_slave_address       : out std_logic_vector(1 downto 0);                     -- address
			switch_pi_avalon_parallel_port_slave_write         : out std_logic;                                        -- write
			switch_pi_avalon_parallel_port_slave_read          : out std_logic;                                        -- read
			switch_pi_avalon_parallel_port_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			switch_pi_avalon_parallel_port_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			switch_pi_avalon_parallel_port_slave_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			switch_pi_avalon_parallel_port_slave_chipselect    : out std_logic;                                        -- chipselect
			sysid_control_slave_address                        : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_address                                  : out std_logic_vector(2 downto 0);                     -- address
			uart_0_s1_write                                    : out std_logic;                                        -- write
			uart_0_s1_read                                     : out std_logic;                                        -- read
			uart_0_s1_readdata                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_writedata                                : out std_logic_vector(15 downto 0);                    -- writedata
			uart_0_s1_begintransfer                            : out std_logic;                                        -- begintransfer
			uart_0_s1_chipselect                               : out std_logic                                         -- chipselect
		);
	end component crypto_wallet_mm_interconnect_0;

	component crypto_wallet_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component crypto_wallet_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_data_master_readdata                                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                               : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                               : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                   : std_logic_vector(26 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                                : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                      : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                                     : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                                 : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                            : std_logic_vector(26 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                               : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_chipselect        : std_logic;                     -- mm_interconnect_0:buttons_pi_avalon_parallel_port_slave_chipselect -> buttons_pi:chipselect
	signal mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_readdata          : std_logic_vector(31 downto 0); -- buttons_pi:readdata -> mm_interconnect_0:buttons_pi_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:buttons_pi_avalon_parallel_port_slave_address -> buttons_pi:address
	signal mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_read              : std_logic;                     -- mm_interconnect_0:buttons_pi_avalon_parallel_port_slave_read -> buttons_pi:read
	signal mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:buttons_pi_avalon_parallel_port_slave_byteenable -> buttons_pi:byteenable
	signal mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_write             : std_logic;                     -- mm_interconnect_0:buttons_pi_avalon_parallel_port_slave_write -> buttons_pi:write
	signal mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:buttons_pi_avalon_parallel_port_slave_writedata -> buttons_pi:writedata
	signal mm_interconnect_0_switch_pi_avalon_parallel_port_slave_chipselect         : std_logic;                     -- mm_interconnect_0:switch_pi_avalon_parallel_port_slave_chipselect -> switch_pi:chipselect
	signal mm_interconnect_0_switch_pi_avalon_parallel_port_slave_readdata           : std_logic_vector(31 downto 0); -- switch_pi:readdata -> mm_interconnect_0:switch_pi_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_switch_pi_avalon_parallel_port_slave_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_pi_avalon_parallel_port_slave_address -> switch_pi:address
	signal mm_interconnect_0_switch_pi_avalon_parallel_port_slave_read               : std_logic;                     -- mm_interconnect_0:switch_pi_avalon_parallel_port_slave_read -> switch_pi:read
	signal mm_interconnect_0_switch_pi_avalon_parallel_port_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:switch_pi_avalon_parallel_port_slave_byteenable -> switch_pi:byteenable
	signal mm_interconnect_0_switch_pi_avalon_parallel_port_slave_write              : std_logic;                     -- mm_interconnect_0:switch_pi_avalon_parallel_port_slave_write -> switch_pi:write
	signal mm_interconnect_0_switch_pi_avalon_parallel_port_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:switch_pi_avalon_parallel_port_slave_writedata -> switch_pi:writedata
	signal mm_interconnect_0_led_po_avalon_parallel_port_slave_chipselect            : std_logic;                     -- mm_interconnect_0:led_po_avalon_parallel_port_slave_chipselect -> led_po:chipselect
	signal mm_interconnect_0_led_po_avalon_parallel_port_slave_readdata              : std_logic_vector(31 downto 0); -- led_po:readdata -> mm_interconnect_0:led_po_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_led_po_avalon_parallel_port_slave_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_po_avalon_parallel_port_slave_address -> led_po:address
	signal mm_interconnect_0_led_po_avalon_parallel_port_slave_read                  : std_logic;                     -- mm_interconnect_0:led_po_avalon_parallel_port_slave_read -> led_po:read
	signal mm_interconnect_0_led_po_avalon_parallel_port_slave_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:led_po_avalon_parallel_port_slave_byteenable -> led_po:byteenable
	signal mm_interconnect_0_led_po_avalon_parallel_port_slave_write                 : std_logic;                     -- mm_interconnect_0:led_po_avalon_parallel_port_slave_write -> led_po:write
	signal mm_interconnect_0_led_po_avalon_parallel_port_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_po_avalon_parallel_port_slave_writedata -> led_po:writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                            : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                            : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                         : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                         : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                                : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                               : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect      : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_chipselect -> epcs_flash_controller:chipselect
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata        : std_logic_vector(31 downto 0); -- epcs_flash_controller:readdata -> mm_interconnect_0:epcs_flash_controller_epcs_control_port_readdata
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_address         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_address -> epcs_flash_controller:address
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_read            : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_read -> mm_interconnect_0_epcs_flash_controller_epcs_control_port_read:in
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_write           : std_logic;                     -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_write -> mm_interconnect_0_epcs_flash_controller_epcs_control_port_write:in
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:epcs_flash_controller_epcs_control_port_writedata -> epcs_flash_controller:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                                     : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                       : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                    : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                        : std_logic_vector(23 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                           : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                                  : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                          : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_uart_0_s1_chipselect                                    : std_logic;                     -- mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	signal mm_interconnect_0_uart_0_s1_readdata                                      : std_logic_vector(15 downto 0); -- uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	signal mm_interconnect_0_uart_0_s1_address                                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_0_s1_address -> uart_0:address
	signal mm_interconnect_0_uart_0_s1_read                                          : std_logic;                     -- mm_interconnect_0:uart_0_s1_read -> mm_interconnect_0_uart_0_s1_read:in
	signal mm_interconnect_0_uart_0_s1_begintransfer                                 : std_logic;                     -- mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	signal mm_interconnect_0_uart_0_s1_write                                         : std_logic;                     -- mm_interconnect_0:uart_0_s1_write -> mm_interconnect_0_uart_0_s1_write:in
	signal mm_interconnect_0_uart_0_s1_writedata                                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	signal irq_mapper_receiver0_irq                                                  : std_logic;                     -- uart_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                  : std_logic;                     -- epcs_flash_controller:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                               : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                            : std_logic;                     -- rst_controller:reset_out -> [buttons_pi:reset, irq_mapper:reset, led_po:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, switch_pi:reset]
	signal rst_controller_reset_out_reset_req                                        : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, epcs_flash_controller:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                             : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in1
	signal reset_reset_n_ports_inv                                                   : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_0_epcs_flash_controller_epcs_control_port_read:inv -> epcs_flash_controller:read_n
	signal mm_interconnect_0_epcs_flash_controller_epcs_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_0_epcs_flash_controller_epcs_control_port_write:inv -> epcs_flash_controller:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                                 : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                                : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_uart_0_s1_read_ports_inv                                : std_logic;                     -- mm_interconnect_0_uart_0_s1_read:inv -> uart_0:read_n
	signal mm_interconnect_0_uart_0_s1_write_ports_inv                               : std_logic;                     -- mm_interconnect_0_uart_0_s1_write:inv -> uart_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, epcs_flash_controller:reset_n, sdram:reset_n, sysid:reset_n, uart_0:reset_n]

begin

	buttons_pi : component crypto_wallet_buttons_pi
		port map (
			clk        => clk_clk,                                                            --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                     --                      reset.reset
			address    => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_readdata,   --                           .readdata
			KEY        => buttons_pi_export                                                   --         external_interface.export
		);

	cpu : component crypto_wallet_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	epcs_flash_controller : component crypto_wallet_epcs_flash_controller
		port map (
			clk        => clk_clk,                                                                   --               clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                                  --             reset.reset_n
			reset_req  => rst_controller_reset_out_reset_req,                                        --                  .reset_req
			address    => mm_interconnect_0_epcs_flash_controller_epcs_control_port_address,         -- epcs_control_port.address
			chipselect => mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect,      --                  .chipselect
			read_n     => mm_interconnect_0_epcs_flash_controller_epcs_control_port_read_ports_inv,  --                  .read_n
			readdata   => mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata,        --                  .readdata
			write_n    => mm_interconnect_0_epcs_flash_controller_epcs_control_port_write_ports_inv, --                  .write_n
			writedata  => mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata,       --                  .writedata
			irq        => irq_mapper_receiver1_irq,                                                  --               irq.irq
			dclk       => epcs_dclk,                                                                 --          external.export
			sce        => epcs_sce,                                                                  --                  .export
			sdo        => epcs_sdo,                                                                  --                  .export
			data0      => epcs_data0                                                                 --                  .export
		);

	led_po : component crypto_wallet_led_po
		port map (
			clk        => clk_clk,                                                        --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                 --                      reset.reset
			address    => mm_interconnect_0_led_po_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_led_po_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_led_po_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_led_po_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_led_po_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_led_po_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_led_po_avalon_parallel_port_slave_readdata,   --                           .readdata
			LEDG       => led_po_export                                                   --         external_interface.export
		);

	sdram : component crypto_wallet_sdram
		port map (
			clk            => clk_clk,                                         --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	switch_pi : component crypto_wallet_switch_pi
		port map (
			clk        => clk_clk,                                                           --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                    --                      reset.reset
			address    => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_readdata,   --                           .readdata
			DIP        => switch_pi_export                                                   --         external_interface.export
		);

	sysid : component crypto_wallet_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	uart_0 : component crypto_wallet_uart_0
		port map (
			clk           => clk_clk,                                     --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_0_uart_0_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_0_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_0_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_0_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_0_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_0_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_0_s1_readdata,        --                    .readdata
			rxd           => uart_0_rxd,                                  -- external_connection.export
			txd           => uart_0_txd,                                  --                    .export
			irq           => irq_mapper_receiver0_irq                     --                 irq.irq
		);

	mm_interconnect_0 : component crypto_wallet_mm_interconnect_0
		port map (
			clk_sys_clk_clk                                    => clk_clk,                                                              --                             clk_sys_clk.clk
			cpu_reset_reset_bridge_in_reset_reset              => rst_controller_reset_out_reset,                                       --         cpu_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                            => cpu_data_master_address,                                              --                         cpu_data_master.address
			cpu_data_master_waitrequest                        => cpu_data_master_waitrequest,                                          --                                        .waitrequest
			cpu_data_master_byteenable                         => cpu_data_master_byteenable,                                           --                                        .byteenable
			cpu_data_master_read                               => cpu_data_master_read,                                                 --                                        .read
			cpu_data_master_readdata                           => cpu_data_master_readdata,                                             --                                        .readdata
			cpu_data_master_write                              => cpu_data_master_write,                                                --                                        .write
			cpu_data_master_writedata                          => cpu_data_master_writedata,                                            --                                        .writedata
			cpu_data_master_debugaccess                        => cpu_data_master_debugaccess,                                          --                                        .debugaccess
			cpu_instruction_master_address                     => cpu_instruction_master_address,                                       --                  cpu_instruction_master.address
			cpu_instruction_master_waitrequest                 => cpu_instruction_master_waitrequest,                                   --                                        .waitrequest
			cpu_instruction_master_read                        => cpu_instruction_master_read,                                          --                                        .read
			cpu_instruction_master_readdata                    => cpu_instruction_master_readdata,                                      --                                        .readdata
			buttons_pi_avalon_parallel_port_slave_address      => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_address,      --   buttons_pi_avalon_parallel_port_slave.address
			buttons_pi_avalon_parallel_port_slave_write        => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_write,        --                                        .write
			buttons_pi_avalon_parallel_port_slave_read         => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_read,         --                                        .read
			buttons_pi_avalon_parallel_port_slave_readdata     => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_readdata,     --                                        .readdata
			buttons_pi_avalon_parallel_port_slave_writedata    => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_writedata,    --                                        .writedata
			buttons_pi_avalon_parallel_port_slave_byteenable   => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_byteenable,   --                                        .byteenable
			buttons_pi_avalon_parallel_port_slave_chipselect   => mm_interconnect_0_buttons_pi_avalon_parallel_port_slave_chipselect,   --                                        .chipselect
			cpu_debug_mem_slave_address                        => mm_interconnect_0_cpu_debug_mem_slave_address,                        --                     cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                          => mm_interconnect_0_cpu_debug_mem_slave_write,                          --                                        .write
			cpu_debug_mem_slave_read                           => mm_interconnect_0_cpu_debug_mem_slave_read,                           --                                        .read
			cpu_debug_mem_slave_readdata                       => mm_interconnect_0_cpu_debug_mem_slave_readdata,                       --                                        .readdata
			cpu_debug_mem_slave_writedata                      => mm_interconnect_0_cpu_debug_mem_slave_writedata,                      --                                        .writedata
			cpu_debug_mem_slave_byteenable                     => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                     --                                        .byteenable
			cpu_debug_mem_slave_waitrequest                    => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                    --                                        .waitrequest
			cpu_debug_mem_slave_debugaccess                    => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                    --                                        .debugaccess
			epcs_flash_controller_epcs_control_port_address    => mm_interconnect_0_epcs_flash_controller_epcs_control_port_address,    -- epcs_flash_controller_epcs_control_port.address
			epcs_flash_controller_epcs_control_port_write      => mm_interconnect_0_epcs_flash_controller_epcs_control_port_write,      --                                        .write
			epcs_flash_controller_epcs_control_port_read       => mm_interconnect_0_epcs_flash_controller_epcs_control_port_read,       --                                        .read
			epcs_flash_controller_epcs_control_port_readdata   => mm_interconnect_0_epcs_flash_controller_epcs_control_port_readdata,   --                                        .readdata
			epcs_flash_controller_epcs_control_port_writedata  => mm_interconnect_0_epcs_flash_controller_epcs_control_port_writedata,  --                                        .writedata
			epcs_flash_controller_epcs_control_port_chipselect => mm_interconnect_0_epcs_flash_controller_epcs_control_port_chipselect, --                                        .chipselect
			led_po_avalon_parallel_port_slave_address          => mm_interconnect_0_led_po_avalon_parallel_port_slave_address,          --       led_po_avalon_parallel_port_slave.address
			led_po_avalon_parallel_port_slave_write            => mm_interconnect_0_led_po_avalon_parallel_port_slave_write,            --                                        .write
			led_po_avalon_parallel_port_slave_read             => mm_interconnect_0_led_po_avalon_parallel_port_slave_read,             --                                        .read
			led_po_avalon_parallel_port_slave_readdata         => mm_interconnect_0_led_po_avalon_parallel_port_slave_readdata,         --                                        .readdata
			led_po_avalon_parallel_port_slave_writedata        => mm_interconnect_0_led_po_avalon_parallel_port_slave_writedata,        --                                        .writedata
			led_po_avalon_parallel_port_slave_byteenable       => mm_interconnect_0_led_po_avalon_parallel_port_slave_byteenable,       --                                        .byteenable
			led_po_avalon_parallel_port_slave_chipselect       => mm_interconnect_0_led_po_avalon_parallel_port_slave_chipselect,       --                                        .chipselect
			sdram_s1_address                                   => mm_interconnect_0_sdram_s1_address,                                   --                                sdram_s1.address
			sdram_s1_write                                     => mm_interconnect_0_sdram_s1_write,                                     --                                        .write
			sdram_s1_read                                      => mm_interconnect_0_sdram_s1_read,                                      --                                        .read
			sdram_s1_readdata                                  => mm_interconnect_0_sdram_s1_readdata,                                  --                                        .readdata
			sdram_s1_writedata                                 => mm_interconnect_0_sdram_s1_writedata,                                 --                                        .writedata
			sdram_s1_byteenable                                => mm_interconnect_0_sdram_s1_byteenable,                                --                                        .byteenable
			sdram_s1_readdatavalid                             => mm_interconnect_0_sdram_s1_readdatavalid,                             --                                        .readdatavalid
			sdram_s1_waitrequest                               => mm_interconnect_0_sdram_s1_waitrequest,                               --                                        .waitrequest
			sdram_s1_chipselect                                => mm_interconnect_0_sdram_s1_chipselect,                                --                                        .chipselect
			switch_pi_avalon_parallel_port_slave_address       => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_address,       --    switch_pi_avalon_parallel_port_slave.address
			switch_pi_avalon_parallel_port_slave_write         => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_write,         --                                        .write
			switch_pi_avalon_parallel_port_slave_read          => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_read,          --                                        .read
			switch_pi_avalon_parallel_port_slave_readdata      => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_readdata,      --                                        .readdata
			switch_pi_avalon_parallel_port_slave_writedata     => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_writedata,     --                                        .writedata
			switch_pi_avalon_parallel_port_slave_byteenable    => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_byteenable,    --                                        .byteenable
			switch_pi_avalon_parallel_port_slave_chipselect    => mm_interconnect_0_switch_pi_avalon_parallel_port_slave_chipselect,    --                                        .chipselect
			sysid_control_slave_address                        => mm_interconnect_0_sysid_control_slave_address,                        --                     sysid_control_slave.address
			sysid_control_slave_readdata                       => mm_interconnect_0_sysid_control_slave_readdata,                       --                                        .readdata
			uart_0_s1_address                                  => mm_interconnect_0_uart_0_s1_address,                                  --                               uart_0_s1.address
			uart_0_s1_write                                    => mm_interconnect_0_uart_0_s1_write,                                    --                                        .write
			uart_0_s1_read                                     => mm_interconnect_0_uart_0_s1_read,                                     --                                        .read
			uart_0_s1_readdata                                 => mm_interconnect_0_uart_0_s1_readdata,                                 --                                        .readdata
			uart_0_s1_writedata                                => mm_interconnect_0_uart_0_s1_writedata,                                --                                        .writedata
			uart_0_s1_begintransfer                            => mm_interconnect_0_uart_0_s1_begintransfer,                            --                                        .begintransfer
			uart_0_s1_chipselect                               => mm_interconnect_0_uart_0_s1_chipselect                                --                                        .chipselect
		);

	irq_mapper : component crypto_wallet_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_epcs_flash_controller_epcs_control_port_read_ports_inv <= not mm_interconnect_0_epcs_flash_controller_epcs_control_port_read;

	mm_interconnect_0_epcs_flash_controller_epcs_control_port_write_ports_inv <= not mm_interconnect_0_epcs_flash_controller_epcs_control_port_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_uart_0_s1_read_ports_inv <= not mm_interconnect_0_uart_0_s1_read;

	mm_interconnect_0_uart_0_s1_write_ports_inv <= not mm_interconnect_0_uart_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of crypto_wallet
